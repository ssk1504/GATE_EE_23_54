
*Title: case(ii) transient analysis

r 1 2 10
V1 1 0 DC 5V
C1 2 0 100u IC=SIN(159*time - PI/4)
.tran 0.002ms 4ms
.control
run
set color0=white
plot v(2)
.endc
.end
