*Title: Case(i)

r 0 1 10
Iin 0 1 SIN(0 1 159)
c 1 0 100u ic=0
.tran 0.02ms 20ms
.control
run
set color0 = white
plot v(1)
.endc
.end
